///////////////////////////////////////////////////////////////////////////////
// Copyright(C) Team . Open source License: MIT.
// ALL RIGHT RESERVED
// File name   : CPU_Defines.svh
// Author      : Juan Jiang
// Date        : 2021-03-20
// Version     : 0.1
// Description :
// none
//    
// Parameter   :没有
//    ...
//    ...
// IO Port     :没有
//    ...
//    ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
//==============================================================================
// 19-06-02 |    Zion    |     0.1     | Original Version
// ...
////////////////////////////////////////////////////////////////////////////////
`ifndef CommonDefines_SVH
`define CommonDefines_SVH

// 这两个定义，感觉大家都能用得到，所以先传上来了。剩下的就等我们都写的差不读之后再一起传上来，现在先各人写各人的
`define WriteEnable 1'b1          // 打开写使能信号
`define WriteDisable 1'b1         // 关闭写使能信号

`endif 