`include "../CommonDefines.svh"
`include "../CPU_Defines.svh"
module ExceptionInEXE(
    input  logic              Overflow_valid,
    input  logic              Trap_valid,
    input  ExceptinPipeType   EXE_ExceptType,
    // 用于产生TLB refetch & 取指令地址错例外
    input  LoadType           EXE_LoadType,
    input  logic              MEM_IsTLBR,
    input  logic              MEM_IsTLBW,
    input  logic [31:0]       MEM_Instr,
    input  logic [4:0]        MEM_Dst,
    input  logic [31:0]       EXE_ALUOut,    // 地址信息

    output ExceptinPipeType   EXE_ExceptType_final
);
// EXE级一共产生5种例外，溢出，trap ，TLBrefetch ， 数据访问地址错误
    assign EXE_ExceptType_final.Interrupt           =  EXE_ExceptType.Interrupt;
    assign EXE_ExceptType_final.WrongAddressinIF    =  EXE_ExceptType.WrongAddressinIF;
    assign EXE_ExceptType_final.ReservedInstruction =  EXE_ExceptType.ReservedInstruction;
    assign EXE_ExceptType_final.CoprocessorUnusable =  EXE_ExceptType.CoprocessorUnusable;
    assign EXE_ExceptType_final.Syscall             =  EXE_ExceptType.Syscall;
    assign EXE_ExceptType_final.Break               =  EXE_ExceptType.Break;
    assign EXE_ExceptType_final.Eret                =  EXE_ExceptType.Eret;
    assign EXE_ExceptType_final.WrWrongAddressinMEM =  EXE_StoreType.DMWr&&(((EXE_StoreType.size == `STORETYPE_SW)&&(EXE_ALUOut[1:0] != 2'b00))||((EXE_StoreType.size == `STORETYPE_SH)&&(EXE_ALUOut[0] != 1'b0)));
    assign EXE_ExceptType_final.RdWrongAddressinMEM =  EXE_LoadType.ReadMem&&(((EXE_LoadType.size == 2'b00)&&(EXE_ALUOut[1:0] != 2'b00))||((EXE_LoadType.size == 2'b01)&&(EXE_ALUOut[0] != 1'b0)));
    assign EXE_ExceptType_final.Overflow            =  Overflow_valid;
    assign EXE_ExceptType_final.TLBRefillinIF       =  EXE_ExceptType.TLBRefillinIF;
    assign EXE_ExceptType_final.TLBInvalidinIF      =  EXE_ExceptType.TLBInvalidinIF;
    assign EXE_ExceptType_final.RdTLBRefillinMEM    =  EXE_ExceptType.RdTLBRefillinMEM;
    assign EXE_ExceptType_final.RdTLBInvalidinMEM   =  EXE_ExceptType.RdTLBInvalidinMEM;
    assign EXE_ExceptType_final.WrTLBRefillinMEM    =  EXE_ExceptType.WrTLBRefillinMEM; 
    assign EXE_ExceptType_final.WrTLBInvalidinMEM   =  EXE_ExceptType.WrTLBInvalidinMEM;   
    assign EXE_ExceptType_final.TLBModified         =  EXE_ExceptType.TLBModified;
    assign EXE_ExceptType_final.Refetch             =  (MEM_IsTLBR == 1'b1 || MEM_IsTLBW == 1'b1 || (MEM_Instr[31:21] == 11'b01000000100 && MEM_Dst == `CP0_REG_ENTRYHI));
    assign EXE_ExceptType_final.Trap                =  Trap_valid;
endmodule