`define WriteEnable 1'b1
`define InterruptNotAssert 1'b0
`define InterruptAssert 1'b1
`define InDelaySlot 1'b1