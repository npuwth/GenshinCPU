/*
 * @Author: your name
 * @Date: 2021-07-06 11:28:11
 * @LastEditTime: 2021-07-06 11:28:14
 * @LastEditors: Please set LastEditors
 * @Description: In User Settings Edit
 * @FilePath: \NewCache\StateMachine.sv
 */
module StateMachine(
    port_list
);
    
endmodule