///////////////////////////////////////////////////////////////////////////////
// Copyright(C) Team . Open source License: MIT.
// ALL RIGHT RESERVED
// File name   : CPU_Defines.svh
// Author      : Juan Jiang
// Date        : 2021-03-20
// Version     : 0.1
// Description :
// none
//    
// Parameter   :没有
//    ...
//    ...
// IO Port     :没有
//    ...
//    ...
// Modification History:
//   Date   |   Author   |   Version   |   Change Description
//==============================================================================
// 19-06-02 |    Zion    |     0.1     | Original Version
// ...
////////////////////////////////////////////////////////////////////////////////
`ifndef CommonDefines_SVH
`define CommonDefines_SVH



`endif CommonDefines_SVH